VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dff
  CLASS BLOCK ;
  FOREIGN dff ;
  ORIGIN 4.650 0.540 ;
  SIZE 22.080 BY 3.760 ;
  PIN D
    ANTENNAGATEAREA 0.253500 ;
    PORT
      LAYER li1 ;
        RECT -2.400 0.720 -1.980 1.080 ;
    END
  END D
  PIN clk
    ANTENNAGATEAREA 0.760500 ;
    PORT
      LAYER li1 ;
        RECT -4.650 1.080 -4.350 1.830 ;
        RECT -0.480 1.530 -0.210 1.800 ;
        RECT 11.430 1.710 11.760 1.770 ;
        RECT 11.250 1.680 11.760 1.710 ;
        RECT 11.010 1.530 11.760 1.680 ;
        RECT -0.570 1.200 -0.150 1.530 ;
        RECT -4.650 0.720 -4.230 1.080 ;
        RECT 2.220 0.810 2.640 1.410 ;
        RECT 11.010 1.320 11.430 1.530 ;
      LAYER met1 ;
        RECT -4.650 1.530 12.000 1.830 ;
        RECT 2.220 1.020 2.640 1.530 ;
    END
  END clk
  PIN Q
    ANTENNADIFFAREA 0.507000 ;
    PORT
      LAYER li1 ;
        RECT 16.800 1.230 17.040 2.440 ;
        RECT 16.860 1.050 17.040 1.230 ;
        RECT 16.860 0.750 17.400 1.050 ;
        RECT 16.860 0.570 17.040 0.750 ;
        RECT 16.800 0.210 17.040 0.570 ;
    END
  END Q
  PIN vss
    ANTENNADIFFAREA 2.028600 ;
    PORT
      LAYER li1 ;
        RECT -4.050 0.210 -3.450 0.570 ;
        RECT -1.800 0.210 -1.200 0.570 ;
        RECT 3.960 0.210 4.560 0.570 ;
        RECT 6.210 0.210 6.810 0.570 ;
        RECT 11.940 0.210 12.540 0.570 ;
        RECT 13.770 0.210 14.370 0.570 ;
        RECT 15.990 0.210 16.590 0.570 ;
        RECT -4.050 -0.120 -3.720 0.210 ;
        RECT -1.800 -0.120 -1.470 0.210 ;
        RECT 3.960 -0.120 4.290 0.210 ;
        RECT 6.210 -0.120 6.540 0.210 ;
        RECT 11.940 -0.120 12.270 0.210 ;
        RECT 13.770 -0.120 14.100 0.210 ;
        RECT 15.990 -0.120 16.320 0.210 ;
      LAYER met1 ;
        RECT -4.290 -0.150 17.310 0.150 ;
    END
  END vss
  PIN vdd
    ANTENNADIFFAREA 6.134100 ;
    PORT
      LAYER nwell ;
        RECT -4.290 1.020 17.250 2.650 ;
      LAYER li1 ;
        RECT -4.050 2.440 -3.720 2.800 ;
        RECT -1.800 2.440 -1.470 2.800 ;
        RECT 3.960 2.440 4.290 2.800 ;
        RECT 6.210 2.440 6.540 2.800 ;
        RECT 11.940 2.440 12.270 2.800 ;
        RECT 13.770 2.440 14.100 2.800 ;
        RECT 15.990 2.440 16.320 2.800 ;
        RECT -4.050 1.230 -3.450 2.440 ;
        RECT -1.800 1.230 -1.200 2.440 ;
        RECT 3.960 1.230 4.560 2.440 ;
        RECT 6.210 1.230 6.810 2.440 ;
        RECT 11.940 1.230 12.540 2.440 ;
        RECT 13.770 1.230 14.370 2.440 ;
        RECT 15.990 1.230 16.590 2.440 ;
      LAYER met1 ;
        RECT -4.290 2.530 17.430 2.830 ;
    END
  END vdd
  OBS
      LAYER li1 ;
        RECT 2.910 2.980 7.260 3.220 ;
        RECT -3.240 0.480 -3.000 2.440 ;
        RECT -0.990 2.230 0.360 2.440 ;
        RECT -3.240 0.270 -2.970 0.480 ;
        RECT -3.240 0.210 -3.000 0.270 ;
        RECT -0.990 0.210 -0.750 2.230 ;
        RECT 0.090 1.230 0.360 2.230 ;
        RECT 0.720 1.200 0.960 2.440 ;
        RECT 1.320 2.020 1.590 2.440 ;
        RECT 2.910 2.020 3.150 2.980 ;
        RECT 1.320 1.770 3.150 2.020 ;
        RECT 1.320 1.230 1.590 1.770 ;
        RECT 0.780 1.020 0.960 1.200 ;
        RECT 0.780 0.840 2.040 1.020 ;
        RECT 0.180 0.720 0.600 0.750 ;
        RECT -0.270 0.420 0.600 0.720 ;
        RECT 1.860 0.600 2.040 0.840 ;
        RECT 1.230 0.210 1.500 0.570 ;
        RECT -0.990 0.030 1.500 0.210 ;
        RECT 1.860 -0.210 2.100 0.600 ;
        RECT 2.460 0.570 2.700 0.600 ;
        RECT 2.460 0.510 2.730 0.570 ;
        RECT 2.940 0.510 3.150 1.770 ;
        RECT 4.770 1.230 5.010 2.440 ;
        RECT 7.020 1.230 7.260 2.980 ;
        RECT 9.300 2.980 15.210 3.220 ;
        RECT 8.070 1.230 8.340 2.440 ;
        RECT 8.700 1.230 8.940 2.440 ;
        RECT 9.300 1.230 9.570 2.980 ;
        RECT 3.360 0.720 3.780 1.080 ;
        RECT 4.830 1.050 5.010 1.230 ;
        RECT 5.610 1.050 6.030 1.080 ;
        RECT 4.830 0.750 6.030 1.050 ;
        RECT 2.460 0.300 3.150 0.510 ;
        RECT 2.460 0.210 2.730 0.300 ;
        RECT 3.450 -0.210 3.720 0.720 ;
        RECT 4.830 0.570 5.010 0.750 ;
        RECT 4.770 0.210 5.010 0.570 ;
        RECT 5.610 0.720 6.030 0.750 ;
        RECT 1.860 -0.450 3.720 -0.210 ;
        RECT 5.610 -0.300 5.880 0.720 ;
        RECT 7.080 0.570 7.260 1.230 ;
        RECT 7.020 0.210 7.260 0.570 ;
        RECT 7.470 0.510 7.890 1.080 ;
        RECT 8.160 -0.300 8.340 1.230 ;
        RECT 8.760 1.050 8.940 1.230 ;
        RECT 8.760 0.870 9.840 1.050 ;
        RECT 9.660 0.570 9.840 0.870 ;
        RECT 10.350 0.570 10.530 2.980 ;
        RECT 12.750 1.230 12.990 2.440 ;
        RECT 14.580 1.230 14.820 2.440 ;
        RECT 10.710 0.720 11.130 1.080 ;
        RECT 11.340 0.720 11.760 1.080 ;
        RECT 12.810 1.050 12.990 1.230 ;
        RECT 13.170 1.050 13.590 1.080 ;
        RECT 12.810 0.750 13.590 1.050 ;
        RECT 9.030 -0.300 9.300 0.570 ;
        RECT 5.610 -0.540 9.300 -0.300 ;
        RECT 9.660 -0.210 9.900 0.570 ;
        RECT 10.260 0.210 10.530 0.570 ;
        RECT 10.770 0.390 11.040 0.720 ;
        RECT 11.340 -0.210 11.580 0.720 ;
        RECT 12.810 0.570 12.990 0.750 ;
        RECT 13.170 0.720 13.590 0.750 ;
        RECT 12.750 0.210 12.990 0.570 ;
        RECT 9.660 -0.450 11.580 -0.210 ;
        RECT 13.410 -0.300 13.590 0.720 ;
        RECT 14.640 1.050 14.820 1.230 ;
        RECT 15.030 1.050 15.210 2.980 ;
        RECT 14.640 0.750 15.210 1.050 ;
        RECT 14.640 0.570 14.820 0.750 ;
        RECT 14.580 0.210 14.820 0.570 ;
        RECT 15.390 0.720 15.810 1.080 ;
        RECT 15.390 -0.300 15.570 0.720 ;
        RECT 13.410 -0.540 15.570 -0.300 ;
      LAYER met1 ;
        RECT 0.180 0.720 0.600 0.750 ;
        RECT -4.320 0.420 12.000 0.720 ;
  END
END dff
END LIBRARY

