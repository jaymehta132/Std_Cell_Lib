magic
tech sky130A
timestamp 1726055963
<< nwell >>
rect -429 102 1725 265
<< nmos >>
rect -342 18 -327 60
rect -117 18 -102 60
rect 153 18 168 60
rect 228 18 243 60
rect 459 18 474 60
rect 684 18 699 60
rect 933 18 948 60
rect 1008 18 1023 60
rect 1257 18 1272 60
rect 1440 18 1455 60
rect 1662 18 1677 60
<< pmos >>
rect -342 120 -327 247
rect -117 120 -102 247
rect 39 120 54 247
rect 114 120 129 247
rect 459 120 474 247
rect 684 120 699 247
rect 837 120 852 247
rect 912 120 927 247
rect 1257 120 1272 247
rect 1440 120 1455 247
rect 1662 120 1677 247
<< ndiff >>
rect -372 48 -342 60
rect -372 30 -366 48
rect -348 30 -342 48
rect -372 18 -342 30
rect -327 48 -297 60
rect -327 30 -321 48
rect -303 30 -297 48
rect -327 18 -297 30
rect -147 48 -117 60
rect -147 30 -141 48
rect -123 30 -117 48
rect -147 18 -117 30
rect -102 48 -72 60
rect -102 30 -96 48
rect -78 30 -72 48
rect 123 48 153 60
rect -102 18 -72 30
rect 123 30 129 48
rect 147 30 153 48
rect 123 18 153 30
rect 168 48 228 60
rect 168 30 189 48
rect 207 30 228 48
rect 168 18 228 30
rect 243 48 273 60
rect 243 30 249 48
rect 267 30 273 48
rect 243 18 273 30
rect 429 48 459 60
rect 429 30 435 48
rect 453 30 459 48
rect 429 18 459 30
rect 474 48 504 60
rect 474 30 480 48
rect 498 30 504 48
rect 474 18 504 30
rect 654 48 684 60
rect 654 30 660 48
rect 678 30 684 48
rect 654 18 684 30
rect 699 48 729 60
rect 699 30 705 48
rect 723 30 729 48
rect 699 18 729 30
rect 903 48 933 60
rect 903 30 909 48
rect 927 30 933 48
rect 903 18 933 30
rect 948 48 1008 60
rect 948 30 969 48
rect 987 30 1008 48
rect 948 18 1008 30
rect 1023 48 1053 60
rect 1023 30 1029 48
rect 1047 30 1053 48
rect 1023 18 1053 30
rect 1227 48 1257 60
rect 1227 30 1233 48
rect 1251 30 1257 48
rect 1227 18 1257 30
rect 1272 48 1302 60
rect 1272 30 1278 48
rect 1296 30 1302 48
rect 1272 18 1302 30
rect 1410 48 1440 60
rect 1410 30 1416 48
rect 1434 30 1440 48
rect 1410 18 1440 30
rect 1455 48 1485 60
rect 1455 30 1461 48
rect 1479 30 1485 48
rect 1455 18 1485 30
rect 1632 48 1662 60
rect 1632 30 1638 48
rect 1656 30 1662 48
rect 1632 18 1662 30
rect 1677 48 1707 60
rect 1677 30 1683 48
rect 1701 30 1707 48
rect 1677 18 1707 30
<< pdiff >>
rect -372 235 -342 247
rect -372 132 -366 235
rect -348 132 -342 235
rect -372 120 -342 132
rect -327 235 -297 247
rect -327 132 -321 235
rect -303 132 -297 235
rect -327 120 -297 132
rect -147 235 -117 247
rect -147 132 -141 235
rect -123 132 -117 235
rect -147 120 -117 132
rect -102 235 -72 247
rect -102 132 -96 235
rect -78 132 -72 235
rect 9 235 39 247
rect -102 120 -72 132
rect 9 132 15 235
rect 33 132 39 235
rect 9 120 39 132
rect 54 235 114 247
rect 54 132 75 235
rect 93 132 114 235
rect 54 120 114 132
rect 129 235 159 247
rect 129 132 135 235
rect 153 132 159 235
rect 129 120 159 132
rect 429 235 459 247
rect 429 132 435 235
rect 453 132 459 235
rect 429 120 459 132
rect 474 235 504 247
rect 474 132 480 235
rect 498 132 504 235
rect 474 120 504 132
rect 654 235 684 247
rect 654 132 660 235
rect 678 132 684 235
rect 654 120 684 132
rect 699 235 729 247
rect 699 132 705 235
rect 723 132 729 235
rect 699 120 729 132
rect 807 235 837 247
rect 807 132 813 235
rect 831 132 837 235
rect 807 120 837 132
rect 852 235 912 247
rect 852 132 873 235
rect 891 132 912 235
rect 852 120 912 132
rect 927 235 957 247
rect 927 132 933 235
rect 951 132 957 235
rect 1227 235 1257 247
rect 927 120 957 132
rect 1227 132 1233 235
rect 1251 132 1257 235
rect 1227 120 1257 132
rect 1272 235 1302 247
rect 1272 132 1278 235
rect 1296 132 1302 235
rect 1272 120 1302 132
rect 1410 235 1440 247
rect 1410 132 1416 235
rect 1434 132 1440 235
rect 1410 120 1440 132
rect 1455 235 1485 247
rect 1455 132 1461 235
rect 1479 132 1485 235
rect 1455 120 1485 132
rect 1632 235 1662 247
rect 1632 132 1638 235
rect 1656 132 1662 235
rect 1632 120 1662 132
rect 1677 235 1707 247
rect 1677 132 1683 235
rect 1701 132 1707 235
rect 1677 120 1707 132
<< ndiffc >>
rect -366 30 -348 48
rect -321 30 -303 48
rect -141 30 -123 48
rect -96 30 -78 48
rect 129 30 147 48
rect 189 30 207 48
rect 249 30 267 48
rect 435 30 453 48
rect 480 30 498 48
rect 660 30 678 48
rect 705 30 723 48
rect 909 30 927 48
rect 969 30 987 48
rect 1029 30 1047 48
rect 1233 30 1251 48
rect 1278 30 1296 48
rect 1416 30 1434 48
rect 1461 30 1479 48
rect 1638 30 1656 48
rect 1683 30 1701 48
<< pdiffc >>
rect -366 132 -348 235
rect -321 132 -303 235
rect -141 132 -123 235
rect -96 132 -78 235
rect 15 132 33 235
rect 75 132 93 235
rect 135 132 153 235
rect 435 132 453 235
rect 480 132 498 235
rect 660 132 678 235
rect 705 132 723 235
rect 813 132 831 235
rect 873 132 891 235
rect 933 132 951 235
rect 1233 132 1251 235
rect 1278 132 1296 235
rect 1416 132 1434 235
rect 1461 132 1479 235
rect 1638 132 1656 235
rect 1683 132 1701 235
<< psubdiff >>
rect -411 48 -372 60
rect -411 30 -402 48
rect -384 30 -372 48
rect -411 18 -372 30
rect -186 48 -147 60
rect -186 30 -177 48
rect -159 30 -147 48
rect -186 18 -147 30
rect 390 48 429 60
rect 390 30 399 48
rect 417 30 429 48
rect 390 18 429 30
rect 615 48 654 60
rect 615 30 624 48
rect 642 30 654 48
rect 615 18 654 30
rect 1188 48 1227 60
rect 1188 30 1197 48
rect 1215 30 1227 48
rect 1188 18 1227 30
rect 1371 48 1410 60
rect 1371 30 1380 48
rect 1398 30 1410 48
rect 1371 18 1410 30
rect 1593 48 1632 60
rect 1593 30 1602 48
rect 1620 30 1632 48
rect 1593 18 1632 30
<< nsubdiff >>
rect -411 235 -372 247
rect -411 132 -402 235
rect -384 132 -372 235
rect -411 120 -372 132
rect -186 235 -147 247
rect -186 132 -177 235
rect -159 132 -147 235
rect -186 120 -147 132
rect 390 235 429 247
rect 390 132 399 235
rect 417 132 429 235
rect 390 120 429 132
rect 615 235 654 247
rect 615 132 624 235
rect 642 132 654 235
rect 615 120 654 132
rect 1188 235 1227 247
rect 1188 132 1197 235
rect 1215 132 1227 235
rect 1188 120 1227 132
rect 1371 235 1410 247
rect 1371 132 1380 235
rect 1398 132 1410 235
rect 1371 120 1410 132
rect 1593 235 1632 247
rect 1593 132 1602 235
rect 1620 132 1632 235
rect 1593 120 1632 132
<< psubdiffcont >>
rect -402 30 -384 48
rect -177 30 -159 48
rect 399 30 417 48
rect 624 30 642 48
rect 1197 30 1215 48
rect 1380 30 1398 48
rect 1602 30 1620 48
<< nsubdiffcont >>
rect -402 132 -384 235
rect -177 132 -159 235
rect 399 132 417 235
rect 624 132 642 235
rect 1197 132 1215 235
rect 1380 132 1398 235
rect 1602 132 1620 235
<< poly >>
rect -342 247 -327 262
rect -117 247 -102 262
rect 39 247 54 262
rect 114 247 129 262
rect 459 247 474 262
rect 684 247 699 262
rect 837 247 852 262
rect 912 247 927 262
rect 1257 247 1272 262
rect 1440 247 1455 262
rect 1662 247 1677 262
rect -57 144 -15 153
rect -57 126 -45 144
rect -27 126 -15 144
rect -57 120 -15 126
rect 1101 159 1143 168
rect 966 141 1113 159
rect 1131 141 1143 159
rect 966 132 1143 141
rect -465 105 -411 108
rect -342 105 -327 120
rect -465 99 -327 105
rect -465 81 -453 99
rect -435 81 -327 99
rect -465 75 -327 81
rect -465 72 -411 75
rect -342 60 -327 75
rect -240 105 -186 108
rect -117 105 -102 120
rect -240 99 -102 105
rect -240 81 -228 99
rect -210 81 -102 99
rect -45 111 -15 120
rect 39 111 54 120
rect -45 96 54 111
rect 114 90 129 120
rect 222 108 264 114
rect 222 90 234 108
rect 252 90 264 108
rect -240 75 -102 81
rect 78 75 168 90
rect 222 78 264 90
rect 336 105 390 108
rect 459 105 474 120
rect 336 99 474 105
rect 336 81 348 99
rect 366 81 474 99
rect -240 72 -186 75
rect -117 60 -102 75
rect 18 69 93 75
rect 18 51 30 69
rect 48 54 93 69
rect 153 60 168 75
rect 228 60 243 78
rect 336 75 474 81
rect 336 72 390 75
rect 459 60 474 75
rect 561 105 615 108
rect 684 105 699 120
rect 837 111 852 120
rect 561 99 699 105
rect 561 81 573 99
rect 591 81 699 99
rect 561 75 699 81
rect 561 72 615 75
rect 684 60 699 75
rect 747 99 852 111
rect 747 81 759 99
rect 777 96 852 99
rect 912 105 927 120
rect 966 105 984 132
rect 777 81 801 96
rect 912 87 984 105
rect 1056 99 1113 108
rect 747 72 801 81
rect 933 60 948 87
rect 1056 84 1083 99
rect 1008 81 1083 84
rect 1101 81 1113 99
rect 1008 72 1113 81
rect 1134 105 1188 108
rect 1257 105 1272 120
rect 1134 99 1272 105
rect 1134 81 1146 99
rect 1164 81 1272 99
rect 1134 75 1272 81
rect 1134 72 1188 75
rect 1008 69 1071 72
rect 1008 60 1023 69
rect 1257 60 1272 75
rect 1317 105 1371 108
rect 1440 105 1455 120
rect 1317 99 1455 105
rect 1317 81 1329 99
rect 1347 81 1455 99
rect 1317 75 1455 81
rect 1317 72 1371 75
rect 1440 60 1455 75
rect 1539 105 1593 108
rect 1662 105 1677 120
rect 1539 99 1677 105
rect 1539 81 1551 99
rect 1569 81 1677 99
rect 1539 75 1677 81
rect 1539 72 1593 75
rect 1662 60 1677 75
rect 48 51 60 54
rect 18 42 60 51
rect -342 3 -327 18
rect -117 3 -102 18
rect 153 3 168 18
rect 228 3 243 18
rect 459 3 474 18
rect 684 3 699 18
rect 933 3 948 18
rect 1008 3 1023 18
rect 1257 3 1272 18
rect 1440 3 1455 18
rect 1662 3 1677 18
<< polycont >>
rect -45 126 -27 144
rect 1113 141 1131 159
rect -453 81 -435 99
rect -228 81 -210 99
rect 234 90 252 108
rect 348 81 366 99
rect 30 51 48 69
rect 573 81 591 99
rect 759 81 777 99
rect 1083 81 1101 99
rect 1146 81 1164 99
rect 1329 81 1347 99
rect 1551 81 1569 99
<< locali >>
rect 291 298 726 322
rect -405 244 -372 256
rect -180 244 -147 256
rect -405 235 -345 244
rect -465 177 -435 183
rect -465 159 -462 177
rect -438 159 -435 177
rect -465 108 -435 159
rect -405 132 -402 235
rect -384 132 -366 235
rect -348 132 -345 235
rect -405 123 -345 132
rect -324 235 -300 244
rect -324 132 -321 235
rect -303 132 -300 235
rect -465 99 -423 108
rect -465 81 -453 99
rect -435 81 -423 99
rect -465 72 -423 81
rect -324 69 -300 132
rect -180 235 -120 244
rect -180 132 -177 235
rect -159 132 -141 235
rect -123 132 -120 235
rect -180 123 -120 132
rect -99 235 36 244
rect -99 132 -96 235
rect -78 223 15 235
rect -78 132 -75 223
rect -48 177 -21 180
rect -48 156 -45 177
rect -24 156 -21 177
rect -48 153 -21 156
rect -240 99 -198 108
rect -240 81 -228 99
rect -210 81 -198 99
rect -240 72 -198 81
rect -405 48 -345 57
rect -405 30 -402 48
rect -384 30 -366 48
rect -348 30 -345 48
rect -405 21 -345 30
rect -180 48 -120 57
rect -324 30 -321 48
rect -303 30 -297 48
rect -324 27 -297 30
rect -180 30 -177 48
rect -159 30 -141 48
rect -123 30 -120 48
rect -324 21 -300 27
rect -180 21 -120 30
rect -99 48 -75 132
rect -57 144 -15 153
rect -57 126 -45 144
rect -27 126 -15 144
rect -57 120 -15 126
rect 9 132 15 223
rect 33 132 36 235
rect 9 123 36 132
rect 72 235 96 244
rect 72 132 75 235
rect 93 132 96 235
rect 72 120 96 132
rect 132 235 159 244
rect 132 132 135 235
rect 153 202 159 235
rect 291 202 315 298
rect 153 177 315 202
rect 153 132 159 177
rect 132 123 159 132
rect 222 138 264 141
rect 78 102 96 120
rect 222 117 231 138
rect 252 117 264 138
rect 222 108 264 117
rect 78 84 204 102
rect 18 72 60 75
rect -99 30 -96 48
rect -78 30 -75 48
rect -27 69 60 72
rect -27 48 -12 69
rect 9 51 30 69
rect 48 51 60 69
rect 186 60 204 84
rect 222 90 234 108
rect 252 90 264 108
rect 222 81 264 90
rect 9 48 60 51
rect -27 42 60 48
rect 123 48 150 57
rect -99 21 -75 30
rect 123 30 129 48
rect 147 30 150 48
rect 123 21 150 30
rect -405 12 -372 21
rect -180 12 -147 21
rect -99 3 150 21
rect 186 48 210 60
rect 186 30 189 48
rect 207 30 210 48
rect 186 -21 210 30
rect 246 57 270 60
rect 246 51 273 57
rect 294 51 315 177
rect 396 244 429 256
rect 621 244 654 256
rect 396 235 456 244
rect 396 132 399 235
rect 417 132 435 235
rect 453 132 456 235
rect 396 123 456 132
rect 477 235 501 244
rect 477 132 480 235
rect 498 132 501 235
rect 477 123 501 132
rect 621 235 681 244
rect 621 132 624 235
rect 642 132 660 235
rect 678 132 681 235
rect 621 123 681 132
rect 702 235 726 298
rect 930 298 1521 322
rect 702 132 705 235
rect 723 132 726 235
rect 702 123 726 132
rect 807 235 834 244
rect 807 132 813 235
rect 831 132 834 235
rect 807 123 834 132
rect 870 235 894 244
rect 870 132 873 235
rect 891 132 894 235
rect 870 123 894 132
rect 930 235 957 298
rect 930 132 933 235
rect 951 132 957 235
rect 930 123 957 132
rect 336 99 378 108
rect 336 81 348 99
rect 366 81 378 99
rect 336 72 378 81
rect 483 105 501 123
rect 561 105 603 108
rect 483 99 603 105
rect 483 81 573 99
rect 591 81 603 99
rect 483 75 603 81
rect 246 48 315 51
rect 246 30 249 48
rect 267 30 315 48
rect 246 21 273 30
rect 345 -21 372 72
rect 483 57 501 75
rect 396 48 456 57
rect 396 30 399 48
rect 417 30 435 48
rect 453 30 456 48
rect 396 21 456 30
rect 477 48 501 57
rect 477 30 480 48
rect 498 30 501 48
rect 477 21 501 30
rect 561 72 603 75
rect 396 12 429 21
rect 186 -45 372 -21
rect 561 -30 588 72
rect 708 57 726 123
rect 621 48 681 57
rect 621 30 624 48
rect 642 30 660 48
rect 678 30 681 48
rect 621 21 681 30
rect 702 48 726 57
rect 747 99 789 108
rect 747 81 759 99
rect 777 81 789 99
rect 747 69 789 81
rect 747 51 753 69
rect 783 51 789 69
rect 702 30 705 48
rect 723 30 726 48
rect 702 21 726 30
rect 621 12 654 21
rect 816 -30 834 123
rect 876 105 894 123
rect 876 87 984 105
rect 966 57 984 87
rect 1035 57 1053 298
rect 1194 244 1227 256
rect 1377 244 1410 256
rect 1194 235 1254 244
rect 1143 174 1176 177
rect 1143 171 1146 174
rect 1125 168 1146 171
rect 1101 159 1146 168
rect 1101 141 1113 159
rect 1131 156 1146 159
rect 1173 156 1176 174
rect 1131 153 1176 156
rect 1131 141 1143 153
rect 1101 132 1143 141
rect 1194 132 1197 235
rect 1215 132 1233 235
rect 1251 132 1254 235
rect 1194 123 1254 132
rect 1275 235 1299 244
rect 1275 132 1278 235
rect 1296 132 1299 235
rect 1275 123 1299 132
rect 1377 235 1437 244
rect 1377 132 1380 235
rect 1398 132 1416 235
rect 1434 132 1437 235
rect 1377 123 1437 132
rect 1458 235 1482 244
rect 1458 132 1461 235
rect 1479 132 1482 235
rect 1458 123 1482 132
rect 1071 99 1113 108
rect 1071 81 1083 99
rect 1101 81 1113 99
rect 1071 72 1113 81
rect 1134 99 1176 108
rect 1134 81 1146 99
rect 1164 81 1176 99
rect 1134 72 1176 81
rect 1281 105 1299 123
rect 1317 105 1359 108
rect 1281 99 1359 105
rect 1281 81 1329 99
rect 1347 81 1359 99
rect 1281 75 1359 81
rect 903 48 930 57
rect 903 30 909 48
rect 927 30 930 48
rect 903 -30 930 30
rect 561 -54 930 -30
rect 966 48 990 57
rect 966 30 969 48
rect 987 30 990 48
rect 966 -21 990 30
rect 1026 48 1053 57
rect 1026 30 1029 48
rect 1047 30 1053 48
rect 1077 66 1104 72
rect 1077 39 1104 48
rect 1026 21 1053 30
rect 1134 -21 1158 72
rect 1281 57 1299 75
rect 1317 72 1359 75
rect 1194 48 1254 57
rect 1194 30 1197 48
rect 1215 30 1233 48
rect 1251 30 1254 48
rect 1194 21 1254 30
rect 1275 48 1299 57
rect 1275 30 1278 48
rect 1296 30 1299 48
rect 1275 21 1299 30
rect 1194 12 1227 21
rect 966 -45 1158 -21
rect 1341 -30 1359 72
rect 1464 105 1482 123
rect 1503 105 1521 298
rect 1599 244 1632 256
rect 1599 235 1659 244
rect 1599 132 1602 235
rect 1620 132 1638 235
rect 1656 132 1659 235
rect 1599 123 1659 132
rect 1680 235 1704 244
rect 1680 132 1683 235
rect 1701 132 1704 235
rect 1680 123 1704 132
rect 1464 75 1521 105
rect 1539 99 1581 108
rect 1539 81 1551 99
rect 1569 81 1581 99
rect 1464 57 1482 75
rect 1377 48 1437 57
rect 1377 30 1380 48
rect 1398 30 1416 48
rect 1434 30 1437 48
rect 1377 21 1437 30
rect 1458 48 1482 57
rect 1458 30 1461 48
rect 1479 30 1482 48
rect 1458 21 1482 30
rect 1539 72 1581 81
rect 1686 105 1704 123
rect 1686 75 1740 105
rect 1377 12 1410 21
rect 1539 -30 1557 72
rect 1686 57 1704 75
rect 1599 48 1659 57
rect 1599 30 1602 48
rect 1620 30 1638 48
rect 1656 30 1659 48
rect 1599 21 1659 30
rect 1680 48 1704 57
rect 1680 30 1683 48
rect 1701 30 1704 48
rect 1680 21 1704 30
rect 1599 12 1632 21
rect 1341 -54 1557 -30
<< viali >>
rect -405 256 -372 280
rect -180 256 -147 280
rect -462 159 -438 177
rect -45 156 -24 177
rect -324 48 -300 69
rect 231 117 252 138
rect -12 48 9 69
rect -405 -12 -372 12
rect -180 -12 -147 12
rect 396 256 429 280
rect 621 256 654 280
rect 396 -12 429 12
rect 753 51 783 69
rect 621 -12 654 12
rect 1194 256 1227 280
rect 1377 256 1410 280
rect 1146 156 1173 174
rect 1077 48 1104 66
rect 1194 -12 1227 12
rect 1599 256 1632 280
rect 1377 -12 1410 12
rect 1599 -12 1632 12
<< metal1 >>
rect -429 280 1743 283
rect -429 256 -405 280
rect -372 256 -180 280
rect -147 256 396 280
rect 429 256 621 280
rect 654 256 1194 280
rect 1227 256 1377 280
rect 1410 256 1599 280
rect 1632 256 1743 280
rect -429 253 1743 256
rect -465 177 1200 183
rect -465 159 -462 177
rect -438 159 -45 177
rect -465 156 -45 159
rect -24 174 1200 177
rect -24 156 1146 174
rect 1173 156 1200 174
rect -465 153 1200 156
rect 222 138 264 153
rect 222 117 231 138
rect 252 117 264 138
rect 222 102 264 117
rect 18 72 60 75
rect -432 69 1200 72
rect -432 48 -324 69
rect -300 48 -12 69
rect 9 51 753 69
rect 783 66 1200 69
rect 783 51 1077 66
rect 9 48 1077 51
rect 1104 48 1200 66
rect -432 42 1200 48
rect -429 12 1731 15
rect -429 -12 -405 12
rect -372 -12 -180 12
rect -147 -12 396 12
rect 429 -12 621 12
rect 654 -12 1194 12
rect 1227 -12 1377 12
rect 1410 -12 1599 12
rect 1632 -12 1731 12
rect -429 -15 1731 -12
<< labels >>
rlabel locali -240 87 -240 87 1 D
port 1 n
rlabel locali -465 87 -465 87 3 clk
port 2 e
rlabel metal1 -429 -6 -429 -6 1 vss
port 4 n
rlabel metal1 -429 268 -429 268 1 vdd
port 5 n
rlabel locali 1740 87 1740 87 7 Q
port 3 w
<< end >>
