magic
tech sky130A
magscale 1 2
timestamp 1726341943
<< nwell >>
rect -644 380 12 724
<< nmos >>
rect -324 216 -294 300
rect -112 216 -82 300
<< pmos >>
rect -324 422 -294 676
rect -112 422 -82 676
<< ndiff >>
rect -394 272 -324 300
rect -394 238 -384 272
rect -350 238 -324 272
rect -394 216 -324 238
rect -294 276 -236 300
rect -294 242 -282 276
rect -248 242 -236 276
rect -294 216 -236 242
rect -182 272 -112 300
rect -182 238 -172 272
rect -138 238 -112 272
rect -182 216 -112 238
rect -82 276 -24 300
rect -82 242 -70 276
rect -36 242 -24 276
rect -82 216 -24 242
<< pdiff >>
rect -394 642 -324 676
rect -394 606 -370 642
rect -336 606 -324 642
rect -394 568 -324 606
rect -394 532 -370 568
rect -336 532 -324 568
rect -394 494 -324 532
rect -394 458 -370 494
rect -336 458 -324 494
rect -394 422 -324 458
rect -294 642 -236 676
rect -294 606 -282 642
rect -248 606 -236 642
rect -294 568 -236 606
rect -294 532 -282 568
rect -248 532 -236 568
rect -294 494 -236 532
rect -294 458 -282 494
rect -248 458 -236 494
rect -294 422 -236 458
rect -182 642 -112 676
rect -182 606 -158 642
rect -124 606 -112 642
rect -182 568 -112 606
rect -182 532 -158 568
rect -124 532 -112 568
rect -182 494 -112 532
rect -182 458 -158 494
rect -124 458 -112 494
rect -182 422 -112 458
rect -82 642 -24 676
rect -82 606 -70 642
rect -36 606 -24 642
rect -82 568 -24 606
rect -82 532 -70 568
rect -36 532 -24 568
rect -82 494 -24 532
rect -82 458 -70 494
rect -36 458 -24 494
rect -82 422 -24 458
<< ndiffc >>
rect -384 238 -350 272
rect -282 242 -248 276
rect -172 238 -138 272
rect -70 242 -36 276
<< pdiffc >>
rect -370 606 -336 642
rect -370 532 -336 568
rect -370 458 -336 494
rect -282 606 -248 642
rect -282 532 -248 568
rect -282 458 -248 494
rect -158 606 -124 642
rect -158 532 -124 568
rect -158 458 -124 494
rect -70 606 -36 642
rect -70 532 -36 568
rect -70 458 -36 494
<< psubdiff >>
rect -572 274 -488 300
rect -572 238 -548 274
rect -514 238 -488 274
rect -572 216 -488 238
<< nsubdiff >>
rect -572 642 -488 676
rect -572 606 -542 642
rect -508 606 -488 642
rect -572 568 -488 606
rect -572 532 -542 568
rect -508 532 -488 568
rect -572 494 -488 532
rect -572 458 -542 494
rect -508 458 -488 494
rect -572 422 -488 458
<< psubdiffcont >>
rect -548 238 -514 274
<< nsubdiffcont >>
rect -542 606 -508 642
rect -542 532 -508 568
rect -542 458 -508 494
<< poly >>
rect -324 676 -294 721
rect -112 676 -82 721
rect -324 384 -294 422
rect -112 384 -82 422
rect -400 374 -294 384
rect -400 338 -384 374
rect -342 338 -294 374
rect -400 326 -294 338
rect -188 374 -82 384
rect -188 338 -172 374
rect -130 338 -82 374
rect -188 326 -82 338
rect -324 300 -294 326
rect -112 300 -82 326
rect -324 180 -294 216
rect -112 180 -82 216
<< polycont >>
rect -384 338 -342 374
rect -172 338 -130 374
<< locali >>
rect -572 740 -488 746
rect -572 704 -560 740
rect -518 704 -488 740
rect -572 642 -488 704
rect -572 606 -542 642
rect -508 606 -488 642
rect -572 568 -488 606
rect -572 532 -542 568
rect -508 532 -488 568
rect -572 494 -488 532
rect -572 458 -542 494
rect -508 458 -488 494
rect -572 434 -488 458
rect -394 740 -328 746
rect -394 704 -382 740
rect -340 704 -328 740
rect -394 642 -328 704
rect -182 740 -116 746
rect -182 704 -170 740
rect -128 704 -116 740
rect -394 606 -370 642
rect -336 606 -328 642
rect -394 568 -328 606
rect -394 532 -370 568
rect -336 532 -328 568
rect -394 494 -328 532
rect -394 458 -370 494
rect -336 458 -328 494
rect -394 434 -328 458
rect -290 642 -238 658
rect -290 606 -282 642
rect -248 606 -238 642
rect -290 568 -238 606
rect -290 532 -282 568
rect -248 532 -238 568
rect -290 494 -238 532
rect -290 458 -282 494
rect -248 458 -238 494
rect -290 384 -238 458
rect -182 642 -116 704
rect -182 606 -158 642
rect -124 606 -116 642
rect -182 568 -116 606
rect -182 532 -158 568
rect -124 532 -116 568
rect -182 494 -116 532
rect -182 458 -158 494
rect -124 458 -116 494
rect -182 434 -116 458
rect -78 642 -26 658
rect -78 606 -70 642
rect -36 606 -26 642
rect -78 568 -26 606
rect -78 532 -70 568
rect -36 532 -26 568
rect -78 494 -26 532
rect -78 458 -70 494
rect -36 458 -26 494
rect -78 384 -26 458
rect -400 374 -324 384
rect -400 338 -384 374
rect -342 338 -324 374
rect -400 326 -324 338
rect -290 374 -112 384
rect -290 338 -172 374
rect -130 338 -112 374
rect -290 326 -112 338
rect -78 326 12 384
rect -572 274 -488 292
rect -572 238 -548 274
rect -514 238 -488 274
rect -572 196 -488 238
rect -572 158 -554 196
rect -504 158 -488 196
rect -572 148 -488 158
rect -394 272 -334 292
rect -394 238 -384 272
rect -350 238 -334 272
rect -394 192 -334 238
rect -290 276 -238 326
rect -290 242 -282 276
rect -248 242 -238 276
rect -290 216 -238 242
rect -182 272 -122 292
rect -182 238 -172 272
rect -138 238 -122 272
rect -394 156 -384 192
rect -342 156 -334 192
rect -394 148 -334 156
rect -182 192 -122 238
rect -78 276 -26 326
rect -78 242 -70 276
rect -36 242 -26 276
rect -78 216 -26 242
rect -182 156 -172 192
rect -130 156 -122 192
rect -182 148 -122 156
<< viali >>
rect -560 704 -518 740
rect -382 704 -340 740
rect -170 704 -128 740
rect -554 158 -504 196
rect -384 156 -342 192
rect -172 156 -130 192
<< metal1 >>
rect -626 740 12 746
rect -626 704 -560 740
rect -518 704 -382 740
rect -340 704 -170 740
rect -128 704 12 740
rect -626 692 12 704
rect -626 196 12 204
rect -626 158 -554 196
rect -504 192 12 196
rect -504 158 -384 192
rect -626 156 -384 158
rect -342 156 -172 192
rect -130 156 12 192
rect -626 148 12 156
<< labels >>
rlabel metal1 -614 166 -614 166 7 Gnd
port 2 w
rlabel locali -398 344 -398 344 7 A
port 3 w
rlabel metal1 -622 730 -622 730 7 Vdd
port 1 w
rlabel locali -4 354 -4 354 3 Z
port 4 e
<< end >>
