magic
tech sky130A
magscale 1 2
timestamp 1726176300
<< nwell >>
rect -644 382 850 724
rect -644 380 -214 382
<< nmos >>
rect -324 216 -294 300
rect -112 216 -82 300
rect -24 216 6 300
rect 422 216 452 300
rect 510 216 540 300
<< pmos >>
rect -324 422 -294 676
rect -112 422 -82 676
rect -24 422 6 676
rect 176 464 206 596
rect 422 422 452 676
rect 510 422 540 676
rect 710 480 740 612
<< ndiff >>
rect -394 272 -324 300
rect -394 238 -384 272
rect -350 238 -324 272
rect -394 216 -324 238
rect -294 276 -236 300
rect -294 242 -282 276
rect -248 242 -236 276
rect -294 216 -236 242
rect -182 272 -112 300
rect -182 238 -172 272
rect -138 238 -112 272
rect -182 216 -112 238
rect -82 276 -24 300
rect -82 242 -70 276
rect -36 242 -24 276
rect -82 216 -24 242
rect 6 276 76 300
rect 6 242 24 276
rect 58 242 76 276
rect 6 216 76 242
rect 352 272 422 300
rect 352 238 362 272
rect 396 238 422 272
rect 352 216 422 238
rect 452 274 510 300
rect 452 240 464 274
rect 498 240 510 274
rect 452 216 510 240
rect 540 276 610 300
rect 540 242 558 276
rect 592 242 610 276
rect 540 216 610 242
<< pdiff >>
rect -394 642 -324 676
rect -394 606 -370 642
rect -336 606 -324 642
rect -394 568 -324 606
rect -394 532 -370 568
rect -336 532 -324 568
rect -394 494 -324 532
rect -394 458 -370 494
rect -336 458 -324 494
rect -394 422 -324 458
rect -294 642 -236 676
rect -294 606 -282 642
rect -248 606 -236 642
rect -294 568 -236 606
rect -294 532 -282 568
rect -248 532 -236 568
rect -294 494 -236 532
rect -294 458 -282 494
rect -248 458 -236 494
rect -294 422 -236 458
rect -170 642 -112 676
rect -170 606 -158 642
rect -124 606 -112 642
rect -170 568 -112 606
rect -170 532 -158 568
rect -124 532 -112 568
rect -170 494 -112 532
rect -170 458 -158 494
rect -124 458 -112 494
rect -170 422 -112 458
rect -82 642 -24 676
rect -82 606 -70 642
rect -36 606 -24 642
rect -82 568 -24 606
rect -82 532 -70 568
rect -36 532 -24 568
rect -82 494 -24 532
rect -82 458 -70 494
rect -36 458 -24 494
rect -82 422 -24 458
rect 6 642 64 676
rect 6 606 18 642
rect 52 606 64 642
rect 6 568 64 606
rect 364 642 422 676
rect 364 606 376 642
rect 410 606 422 642
rect 6 532 18 568
rect 52 532 64 568
rect 6 494 64 532
rect 6 458 18 494
rect 52 458 64 494
rect 118 550 176 596
rect 118 516 130 550
rect 164 516 176 550
rect 118 464 176 516
rect 206 552 264 596
rect 206 518 218 552
rect 252 518 264 552
rect 206 464 264 518
rect 364 568 422 606
rect 364 532 376 568
rect 410 532 422 568
rect 364 494 422 532
rect 6 422 64 458
rect 364 458 376 494
rect 410 458 422 494
rect 364 422 422 458
rect 452 642 510 676
rect 452 606 464 642
rect 498 606 510 642
rect 452 568 510 606
rect 452 532 464 568
rect 498 532 510 568
rect 452 494 510 532
rect 452 458 464 494
rect 498 458 510 494
rect 452 422 510 458
rect 540 642 598 676
rect 540 606 552 642
rect 586 606 598 642
rect 540 568 598 606
rect 540 532 552 568
rect 586 532 598 568
rect 540 494 598 532
rect 540 458 552 494
rect 586 458 598 494
rect 652 568 710 612
rect 652 532 664 568
rect 698 532 710 568
rect 652 480 710 532
rect 740 568 798 612
rect 740 534 752 568
rect 786 534 798 568
rect 740 480 798 534
rect 540 422 598 458
<< ndiffc >>
rect -384 238 -350 272
rect -282 242 -248 276
rect -172 238 -138 272
rect -70 242 -36 276
rect 24 242 58 276
rect 362 238 396 272
rect 464 240 498 274
rect 558 242 592 276
<< pdiffc >>
rect -370 606 -336 642
rect -370 532 -336 568
rect -370 458 -336 494
rect -282 606 -248 642
rect -282 532 -248 568
rect -282 458 -248 494
rect -158 606 -124 642
rect -158 532 -124 568
rect -158 458 -124 494
rect -70 606 -36 642
rect -70 532 -36 568
rect -70 458 -36 494
rect 18 606 52 642
rect 376 606 410 642
rect 18 532 52 568
rect 18 458 52 494
rect 130 516 164 550
rect 218 518 252 552
rect 376 532 410 568
rect 376 458 410 494
rect 464 606 498 642
rect 464 532 498 568
rect 464 458 498 494
rect 552 606 586 642
rect 552 532 586 568
rect 552 458 586 494
rect 664 532 698 568
rect 752 534 786 568
<< psubdiff >>
rect -572 274 -488 300
rect -572 238 -548 274
rect -514 238 -488 274
rect -572 216 -488 238
<< nsubdiff >>
rect -572 642 -488 676
rect -572 606 -542 642
rect -508 606 -488 642
rect -572 568 -488 606
rect -572 532 -542 568
rect -508 532 -488 568
rect -572 494 -488 532
rect -572 458 -542 494
rect -508 458 -488 494
rect -572 422 -488 458
<< psubdiffcont >>
rect -548 238 -514 274
<< nsubdiffcont >>
rect -542 606 -508 642
rect -542 532 -508 568
rect -542 458 -508 494
<< poly >>
rect -324 676 -294 721
rect -112 676 -82 721
rect -24 676 6 721
rect 176 596 206 721
rect 422 676 452 721
rect 510 676 540 721
rect -324 384 -294 422
rect -112 384 -82 422
rect -24 384 6 422
rect 176 384 206 464
rect 710 612 740 721
rect -400 374 -294 384
rect -400 338 -384 374
rect -342 338 -294 374
rect -400 326 -294 338
rect -188 374 206 384
rect -188 338 -172 374
rect -130 338 206 374
rect -188 326 206 338
rect 422 384 452 422
rect 510 384 540 422
rect 710 384 740 480
rect 422 374 740 384
rect 422 338 454 374
rect 496 338 740 374
rect 422 326 740 338
rect -324 300 -294 326
rect -112 300 -82 326
rect -24 300 6 326
rect 422 300 452 326
rect 510 300 540 326
rect -324 180 -294 216
rect -112 180 -82 216
rect -24 180 6 216
rect 422 180 452 216
rect 510 180 540 216
<< polycont >>
rect -384 338 -342 374
rect -172 338 -130 374
rect 454 338 496 374
<< locali >>
rect -572 740 -488 746
rect -572 704 -560 740
rect -518 704 -488 740
rect -572 642 -488 704
rect -572 606 -542 642
rect -508 606 -488 642
rect -572 568 -488 606
rect -572 532 -542 568
rect -508 532 -488 568
rect -572 494 -488 532
rect -572 458 -542 494
rect -508 458 -488 494
rect -572 434 -488 458
rect -394 740 -328 746
rect -394 704 -382 740
rect -340 704 -328 740
rect -394 642 -328 704
rect 366 736 418 746
rect 366 702 376 736
rect 410 702 418 736
rect -394 606 -370 642
rect -336 606 -328 642
rect -394 568 -328 606
rect -394 532 -370 568
rect -336 532 -328 568
rect -394 494 -328 532
rect -394 458 -370 494
rect -336 458 -328 494
rect -394 434 -328 458
rect -290 642 -238 658
rect -290 606 -282 642
rect -248 606 -238 642
rect -290 568 -238 606
rect -290 532 -282 568
rect -248 532 -238 568
rect -290 494 -238 532
rect -290 458 -282 494
rect -248 458 -238 494
rect -290 384 -238 458
rect -168 642 -116 658
rect -168 606 -158 642
rect -124 606 -116 642
rect -168 568 -116 606
rect -168 532 -158 568
rect -124 532 -116 568
rect -168 494 -116 532
rect -168 458 -158 494
rect -124 458 -116 494
rect -168 434 -116 458
rect -78 642 -26 658
rect -78 606 -70 642
rect -36 606 -26 642
rect -78 568 -26 606
rect -78 532 -70 568
rect -36 532 -26 568
rect -78 494 -26 532
rect -78 458 -70 494
rect -36 458 -26 494
rect -400 374 -324 384
rect -400 338 -384 374
rect -342 338 -324 374
rect -400 326 -324 338
rect -290 374 -112 384
rect -290 338 -172 374
rect -130 338 -112 374
rect -290 326 -112 338
rect -572 274 -488 292
rect -572 238 -548 274
rect -514 238 -488 274
rect -572 196 -488 238
rect -572 158 -554 196
rect -504 158 -488 196
rect -572 148 -488 158
rect -394 272 -334 292
rect -394 238 -384 272
rect -350 238 -334 272
rect -394 192 -334 238
rect -290 276 -238 326
rect -290 242 -282 276
rect -248 242 -238 276
rect -290 216 -238 242
rect -182 272 -124 292
rect -182 238 -172 272
rect -138 238 -124 272
rect -394 156 -384 192
rect -342 156 -334 192
rect -394 148 -334 156
rect -182 196 -124 238
rect -78 276 -26 458
rect 10 642 62 658
rect 10 606 18 642
rect 52 606 62 642
rect 10 568 62 606
rect 366 642 418 702
rect 544 736 596 746
rect 544 702 552 736
rect 586 702 596 736
rect 366 606 376 642
rect 410 606 418 642
rect 10 532 18 568
rect 52 532 62 568
rect 10 494 62 532
rect 10 458 18 494
rect 52 458 62 494
rect 120 550 172 596
rect 120 516 130 550
rect 164 516 172 550
rect 120 476 172 516
rect 208 552 260 596
rect 208 518 218 552
rect 252 518 260 552
rect 10 434 62 458
rect -78 242 -70 276
rect -36 242 -26 276
rect -78 216 -26 242
rect 8 276 76 292
rect 8 242 24 276
rect 58 242 76 276
rect -182 158 -170 196
rect -132 158 -124 196
rect -182 148 -124 158
rect 8 196 76 242
rect 208 276 260 518
rect 366 568 418 606
rect 366 532 376 568
rect 410 532 418 568
rect 366 494 418 532
rect 366 458 376 494
rect 410 458 418 494
rect 366 434 418 458
rect 456 642 508 658
rect 456 606 464 642
rect 498 606 508 642
rect 456 568 508 606
rect 456 532 464 568
rect 498 532 508 568
rect 456 494 508 532
rect 456 458 464 494
rect 498 458 508 494
rect 456 434 508 458
rect 544 642 596 702
rect 544 606 552 642
rect 586 606 596 642
rect 742 736 794 746
rect 742 702 750 736
rect 784 702 794 736
rect 544 568 596 606
rect 544 532 552 568
rect 586 532 596 568
rect 544 494 596 532
rect 544 458 552 494
rect 586 458 596 494
rect 654 568 706 612
rect 654 532 664 568
rect 698 532 706 568
rect 654 492 706 532
rect 742 568 794 702
rect 742 534 752 568
rect 786 534 794 568
rect 742 492 794 534
rect 544 434 596 458
rect 438 374 514 384
rect 438 338 454 374
rect 496 338 514 374
rect 438 326 514 338
rect 208 242 218 276
rect 252 242 260 276
rect 208 236 260 242
rect 352 272 410 292
rect 352 238 362 272
rect 396 238 410 272
rect 8 158 14 196
rect 52 158 76 196
rect 8 148 76 158
rect 352 196 410 238
rect 456 274 508 292
rect 456 240 464 274
rect 498 240 508 274
rect 456 216 508 240
rect 542 276 610 292
rect 542 242 558 276
rect 592 242 610 276
rect 352 158 364 196
rect 402 158 410 196
rect 352 148 410 158
rect 542 196 610 242
rect 542 158 548 196
rect 586 158 610 196
rect 542 148 610 158
<< viali >>
rect -560 704 -518 740
rect -382 704 -340 740
rect 376 702 410 736
rect -158 606 -124 642
rect -158 532 -124 568
rect -158 458 -124 494
rect -554 158 -504 196
rect -384 156 -342 192
rect 18 606 52 642
rect 552 702 586 736
rect 18 532 52 568
rect 18 458 52 494
rect 130 516 164 550
rect -70 242 -36 276
rect -170 158 -132 196
rect 464 606 498 642
rect 464 532 498 568
rect 464 458 498 494
rect 750 702 784 736
rect 664 532 698 568
rect 218 242 252 276
rect 14 158 52 196
rect 464 240 498 274
rect 364 158 402 196
rect 548 158 586 196
<< metal1 >>
rect -626 740 850 746
rect -626 704 -560 740
rect -518 704 -382 740
rect -340 736 850 740
rect -340 704 376 736
rect -626 702 376 704
rect 410 702 552 736
rect 586 702 750 736
rect 784 702 850 736
rect -626 692 850 702
rect -170 642 708 658
rect -170 606 -158 642
rect -124 606 18 642
rect 52 606 464 642
rect 498 606 708 642
rect -170 568 708 606
rect -170 532 -158 568
rect -124 532 18 568
rect 52 550 464 568
rect 52 532 130 550
rect -170 516 130 532
rect 164 532 464 550
rect 498 532 664 568
rect 698 532 708 568
rect 164 516 708 532
rect -170 494 708 516
rect -170 458 -158 494
rect -124 458 18 494
rect 52 458 464 494
rect 498 458 708 494
rect -170 434 708 458
rect -82 276 510 282
rect -82 242 -70 276
rect -36 242 218 276
rect 252 274 510 276
rect 252 242 464 274
rect -82 240 464 242
rect 498 240 510 274
rect -82 234 510 240
rect -626 196 850 204
rect -626 158 -554 196
rect -504 192 -170 196
rect -504 158 -384 192
rect -626 156 -384 158
rect -342 158 -170 192
rect -132 158 14 196
rect 52 158 364 196
rect 402 158 548 196
rect 586 158 850 196
rect -342 156 850 158
rect -626 148 850 156
<< labels >>
rlabel metal1 12 736 12 736 1 vdd
port 4 n
rlabel locali 10 174 10 174 1 vss
port 5 n
rlabel locali 444 350 444 350 1 B
port 2 n
rlabel metal1 304 256 304 256 1 Y
port 3 n
rlabel locali -396 346 -396 346 1 A
port 1 n
<< end >>
